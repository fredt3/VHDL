LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY LOCKBRAIN IS
PORT(

KEYPAD	: IN STD_LOGIC_VECTOR (3 DOWNTO 0); 
CLOCK		: IN STD_LOGIC;
ENTER		: IN STD_LOGIC;
RESET		: IN STD_LOGIC;

LED		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0) --MSB is Green LED
);
END LOCKBRAIN;

ARCHITECTURE ARCH OF LOCKBRAIN IS

TYPE state_type IS (
						KEY3, KEY2, KEY1, KEY0, WAITING_KEY3, WAITING_KEY2, WAITING_KEY1, WAITING_KEY0,
						READ_KEY3, READ_KEY2, READ_KEY1, READ_KEY0, TRY13, TRY12, TRY11, TRY10, TRY23,
						TRY22, TRY21, TRY20, TRY33, TRY32, TRY31, TRY30, WAITING_TRY13, WAITING_TRY12,
						WAITING_TRY11, WAITING_TRY10, WAITING_TRY23, WAITING_TRY22, WAITING_TRY21,
						WAITING_TRY20,	WAITING_TRY33, WAITING_TRY32, WAITING_TRY31, WAITING_TRY30, 
						READ_TRY13, READ_TRY12,	READ_TRY11, READ_TRY10, READ_TRY23, READ_TRY22, READ_TRY21,
						READ_TRY20, READ_TRY33,	READ_TRY32, READ_TRY31, READ_TRY30, LOCKED, OPENED);
SIGNAL pr_state, nx_state : state_type := KEY3;
SIGNAL PASSWORD : STD_LOGIC_VECTOR (15 DOWNTO 0);
SIGNAL ATTEMPT : STD_LOGIC_VECTOR (15 DOWNTO 0);
SIGNAL PASSWORD_3, PASSWORD_2, PASSWORD_1, PASSWORD_0 : STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL TRY_3, TRY_2, TRY_1, TRY_0 : STD_LOGIC_VECTOR (3 DOWNTO 0);

BEGIN

PROCESS (PASSWORD_3, PASSWORD_2, PASSWORD_1, PASSWORD_0, TRY_3, TRY_2, TRY_1, TRY_0)
BEGIN --add all the keys together into one password/attempt
	PASSWORD <= PASSWORD_3 & PASSWORD_2 & PASSWORD_1 & PASSWORD_0;
	ATTEMPT <= TRY_3 & TRY_2 & TRY_1 & TRY_0;
END PROCESS;

PROCESS (RESET, CLOCK) --starts program back to creating the password
BEGIN 
	IF (RESET = '0') THEN
		PR_STATE <= KEY3;
	ELSIF (CLOCK'EVENT AND CLOCK = '1') THEN
		PR_STATE <= NX_STATE;
	END IF;
END PROCESS;

PROCESS(PR_STATE, CLOCK, KEYPAD)
BEGIN
CASE PR_STATE IS
--CREATE PASSWORD
WHEN KEY3 =>
	IF (KEYPAD = "1111") THEN --nothing is being pressed
		NX_STATE <= KEY3;
	ELSE								--sees pressing so moves on to next state
		NX_STATE <= READ_KEY3;
	END IF;
	LED <= "1111";					--all lights on to show that you are creating the password
WHEN READ_KEY3 =>
		PASSWORD_3 <= KEYPAD;
		NX_STATE <= WAITING_KEY3;
	LED <= "1111";

WHEN WAITING_KEY3 =>				--checks when you are done pressing the key
	IF (KEYPAD = "1111") THEN
			NX_STATE <= KEY2;
	ELSE
		NX_STATE <= WAITING_KEY3;
	END IF;
	LED <= "1111";
	
WHEN KEY2 =>						--repeats above except now with the 2 number in the password
	IF (KEYPAD = "1111") THEN
		NX_STATE <= KEY2;
	ELSE
		NX_STATE <= READ_KEY2;
	END IF;
	LED <= "1111";
WHEN READ_KEY2 =>
		PASSWORD_2 <= KEYPAD;
		NX_STATE <= WAITING_KEY2;
		LED <= "1111";

WHEN WAITING_KEY2 =>
	IF (KEYPAD = "1111") THEN
		NX_STATE <= KEY1;
	ELSE
		NX_STATE <= WAITING_KEY2;
	END IF;
	LED <= "1111";
	
WHEN KEY1 =>		--third number
	IF (KEYPAD = "1111") THEN
		NX_STATE <= KEY1;
	ELSE
		NX_STATE <= READ_KEY1;
	END IF;
	LED <= "1111";
WHEN READ_KEY1 =>
		PASSWORD_1 <= KEYPAD;
		NX_STATE <= WAITING_KEY1;
		LED <= "1111";

WHEN WAITING_KEY1 =>
	IF (KEYPAD = "1111") THEN
		NX_STATE <= KEY0;
	ELSE
		NX_STATE <= WAITING_KEY1;
	END IF;
	LED <= "1111";
	
WHEN KEY0 =>  --last number
	IF (KEYPAD = "1111") THEN
		NX_STATE <= KEY0;
	ELSE
		NX_STATE <= READ_KEY0;
	END IF;
	LED <= "1111";
WHEN READ_KEY0 =>
		PASSWORD_0 <= KEYPAD;
		NX_STATE <= WAITING_KEY0;
		LED <= "1111";

WHEN WAITING_KEY0 =>
	IF (KEYPAD = "1111") THEN
			IF (ENTER = '0') THEN --stays in this state until enter is pressed, goes onto the attempt
				NX_STATE <= TRY13;
			ELSE
				NX_STATE <= WAITING_KEY0;
			END IF;
	ELSE
		NX_STATE <= WAITING_KEY0;
	END IF;
	LED <= "1111";
	
--ATTEMPT 1	
WHEN TRY13 => --same setup with creating password but with attempting
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY13;
	ELSE
		NX_STATE <= READ_TRY13;
	END IF;
		LED <= "0000"; --no wrong attempts
	
WHEN READ_TRY13 =>
		TRY_3 <= KEYPAD;
		NX_STATE <= WAITING_TRY13;
		LED <= "0000";
	
WHEN WAITING_TRY13 =>
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY12;
	ELSE
		NX_STATE <= WAITING_TRY13;
	END IF;
		LED <= "0000";
	
WHEN TRY12 => --1st attempt 2nd number
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY12;
	ELSE
		NX_STATE <= READ_TRY12;
	END IF;
		LED <= "0000";
	
WHEN READ_TRY12 =>
		TRY_2 <= KEYPAD;
		NX_STATE <= WAITING_TRY12;
		LED <= "0000";
	
WHEN WAITING_TRY12 =>
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY11;
	ELSE
		NX_STATE <= WAITING_TRY12;
	END IF;
		LED <= "0000";

WHEN TRY11 => --1st attempt 3rd number
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY11;
	ELSE
		NX_STATE <= READ_TRY11;
	END IF;
		LED <= "0000";
	
WHEN READ_TRY11 =>
		TRY_1 <= KEYPAD;
		NX_STATE <= WAITING_TRY11;
		LED <= "0000";
	
WHEN WAITING_TRY11 =>
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY10;
	ELSE
		NX_STATE <= WAITING_TRY11;
	END IF;
		LED <= "0000";

WHEN TRY10 => --1st attempt 4th number
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY10;
	ELSE
		NX_STATE <= READ_TRY10;
	END IF;
		LED <= "0000";
	
WHEN READ_TRY10 =>
		TRY_0 <= KEYPAD;
		NX_STATE <= WAITING_TRY10;
		LED <= "0000";
	
WHEN WAITING_TRY10 =>
	IF (KEYPAD = "1111") THEN
			IF (ENTER = '0') THEN
				IF (PASSWORD = ATTEMPT) THEN --sees if attempt is the same as the password
					NX_STATE <= OPENED;
				ELSE
					NX_STATE <= TRY23;
				END IF;
			ELSE
				NX_STATE <= WAITING_TRY10;
			END IF;
	ELSE
		NX_STATE <= WAITING_TRY10;
	END IF;
	LED <= "0000";
	
--ATTEMPT 2
WHEN TRY23 => --same as attempt 1
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY23;
	ELSE
		NX_STATE <= READ_TRY23;
	END IF;
		LED <= "0001"; --one wrong attempt so far
	
WHEN READ_TRY23 =>
		TRY_3 <= KEYPAD;
		NX_STATE <= WAITING_TRY23;
		LED <= "0001";
	
WHEN WAITING_TRY23 =>
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY22;
	ELSE
		NX_STATE <= WAITING_TRY23;
	END IF;
		LED <= "0001";
	
WHEN TRY22 =>
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY22;
	ELSE
		NX_STATE <= READ_TRY22;
	END IF;
		LED <= "0001";
	
WHEN READ_TRY22 =>
		TRY_2 <= KEYPAD;
		NX_STATE <= WAITING_TRY22;
		LED <= "0001";
	
WHEN WAITING_TRY22 =>
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY21;
	ELSE
		NX_STATE <= WAITING_TRY22;
	END IF;
		LED <= "0001";

WHEN TRY21 =>
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY21;
	ELSE
		NX_STATE <= READ_TRY21;
	END IF;
		LED <= "0001";
	
WHEN READ_TRY21 =>
		TRY_1 <= KEYPAD;
		NX_STATE <= WAITING_TRY21;
		LED <= "0001";
	
WHEN WAITING_TRY21 =>
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY20;
	ELSE
		NX_STATE <= WAITING_TRY21;
	END IF;
		LED <= "0001";

WHEN TRY20 =>
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY20;
	ELSE
		NX_STATE <= READ_TRY20;
	END IF;
		LED <= "0001";
	
WHEN READ_TRY20 =>
		TRY_0 <= KEYPAD;
		NX_STATE <= WAITING_TRY20;
		LED <= "0001";
	
WHEN WAITING_TRY20 =>
	IF (KEYPAD = "1111") THEN
			IF (ENTER = '0') THEN
				IF (PASSWORD = ATTEMPT) THEN
					NX_STATE <= OPENED;
				ELSE
					NX_STATE <= TRY33;
				END IF;
			ELSE
				NX_STATE <= WAITING_TRY20;
			END IF;
	ELSE
		NX_STATE <= WAITING_TRY20;
	END IF;
	LED <= "0001";

--ATTEMPT 3
WHEN TRY33 =>
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY33;
	ELSE
		NX_STATE <= READ_TRY33;
	END IF;
		LED <= "0011"; --2 wrong attempts so far
	
WHEN READ_TRY33 =>
		TRY_3 <= KEYPAD;
		NX_STATE <= WAITING_TRY33;
		LED <= "0011";
	
WHEN WAITING_TRY33 =>
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY32;
	ELSE
		NX_STATE <= WAITING_TRY33;
	END IF;
		LED <= "0011";
	
WHEN TRY32 =>
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY32;
	ELSE
		NX_STATE <= READ_TRY32;
	END IF;
		LED <= "0011";
	
WHEN READ_TRY32 =>
		TRY_2 <= KEYPAD;
		NX_STATE <= WAITING_TRY32;
		LED <= "0011";
	
WHEN WAITING_TRY32 =>
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY31;
	ELSE
		NX_STATE <= WAITING_TRY32;
	END IF;
		LED <= "0011";

WHEN TRY31 =>
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY31;
	ELSE
		NX_STATE <= READ_TRY31;
	END IF;
		LED <= "0011";
	
WHEN READ_TRY31 =>
		TRY_1 <= KEYPAD;
		NX_STATE <= WAITING_TRY31;
		LED <= "0011";
	
WHEN WAITING_TRY31 =>
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY30;
	ELSE
		NX_STATE <= WAITING_TRY31;
	END IF;
		LED <= "0011";

WHEN TRY30 =>
	IF (KEYPAD = "1111") THEN
		NX_STATE <= TRY30;
	ELSE
		NX_STATE <= READ_TRY30;
	END IF;
		LED <= "0011";
	
WHEN READ_TRY30 =>
		TRY_0 <= KEYPAD;
		NX_STATE <= WAITING_TRY30;
		LED <= "0011";
	
WHEN WAITING_TRY30 =>
	IF (KEYPAD = "1111") THEN
			IF (ENTER = '0') THEN
				IF (PASSWORD = ATTEMPT) THEN
					NX_STATE <= OPENED;
				ELSE
					NX_STATE <= LOCKED; --not correct locks forever
				END IF;
			ELSE
				NX_STATE <= WAITING_TRY30;
			END IF;
	ELSE
		NX_STATE <= WAITING_TRY30;
	END IF;
	LED <= "0011";	
	
WHEN LOCKED =>
	NX_STATE <= LOCKED;
	LED <= "0111"; --three wrong attempts
	
WHEN OPENED =>
	NX_STATE <= OPENED;
	LED <= "1000"; --correct
	
END CASE;
END PROCESS;
END arch;